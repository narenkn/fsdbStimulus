

module Rxor(output bit [7:0] y, output bit [7:0]  a, output bit [7:0] b, output bit [7:0] count);

endmodule // xor
